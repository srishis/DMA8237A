module dmaTimingControl(dma_if.DUT dif, dmaControlIf cif, dmaRegIf.FSM rif);

import DmaPackage::*; 

// Initial state condition
always_ff @(posedge dif.CLK) state <= SI;
else		             state <= nextstate;
   
// Program condition
always_comb begin
if(IDLE_CYCLE && !dif.CS_N && !dif.HLDA) cif.Program = 1; 
else if(ACTIVE_CYCLE)			 cif.Program = 0;
end

// Write extend
always_comb begin
if(cif.checkWriteExtend)
	if (rif.commandReg[5] == 1'b1 && rif.modeReg[0][3:2] == 2'b01 || rif.modeReg[1][3:2] == 2'b01 || rif.modeReg[2][3:2] == 2'b01 || rif.modeReg[3][3:2] == 2'b01)
	       cif.writeExtend = 1'b1; //fsm read and extended write next state
	else   cif.writeExtend = 1'b0;
else	       cif.writeExtend = 1'b0;
end

// Read or Write operation
always_comb begin
if(cif.checkReadWrite)
	if(rif.modeReg[3:2] == 2'b01 && rif.commandReg[0] == 1'b0 && rif.commandReg[5] == 1'b1) cif.iow = 1'b0;    
	else if(rif.modeReg[3:2] == 2'b10 && rif.commandReg[0] == 1'b0)    			cif.ior = 1'b0;    
else    begin cif.iow = 1'b1; cif.ior = 1'b1; end
end

// End of process by terminal count 
always_comb begin
if(cif.checkEOP )
	if(rif.statusReg[3:0]) cif.eop = 1'b0;  
	else		       cif.eop = 1'b1;
else			       cif.eop = 1'b1;

// Next state logic
always_comb begin   

        nextstate = state;      //default value for nextstate
              
        unique case(1'b1)       // reverse case       
            state[iSI] :
			begin
			if(VALID_DREQ0 || VALID_DREQ1 || VALID_DREQ2 || VALID_DREQ3) 	nextstate = S0;
			else  								nextstate = SI;
			end
			 
            state[iS0] :
			begin
			if(dif.HLDA) 							nextstate = S1;
			else if(!dif.HLDA) 						nextstate = S0;
			else if(!dif.EOP_N) 						nextstate = SI;
			end
			
            state[iS1] :
			begin
			if(!dif.EOP_N) 						        nextstate = SI;
			else								nextstate = S2;
			end
			
            state[iS2] :  
                        begin
			if(!dif.EOP_N) 						        nextstate = SI;
                        else if(!cif.writeExtend)                                       nextstate = S4;   //if write extension not set next state will be S4 
			else if(cif.writeExtend)					nextstate = S3;
                        end

            state[iS3] :
                        begin
			if(!dif.EOP_N) 						        nextstate = SI;
			else								nextstate = S4;
                        end 
			
            state[iS4] :								nextstate = SI;
 
														
        endcase
end
	  
// Output logic
always_comb begin 

// default values for control outputs
{cif.aen, cif.adstb, cif.Program, ACTIVE_CYCLE, IDLE_CYCLE, cif.checkEOP, cif.checkReadWrite, cif.checkWriteExtend} = 8'b00000000;  
{cif.ldCurrAddrTemp, cif.ldCurrWordTemp, cif.ldtempCurrAddr, cif.ldtempCurrWord, cif.enCurrAddr, cif.enCurrWord, } = 6'b000000; 
{cif.validDACK,  cif.writeExtend} = 2'b00;    		 

    unique case(1'b1)  // reverse case

	    state[iSI]: begin IDLE_CYCLE = 1'b1; cif.hrq = 1'b1;  end

	    state[iS0]: begin ACTIVE_CYCLE = 1'b1; cif.hrq = 1'b1; end
				
	    state[iS1]: begin cif.aen = 1'b1; cif.adstb = 1'b1; cif.validDACK = 1'b1; cif.enCurrAddr = 1'b1; cif.enCurrWord = 1'b1; cif.ldCurrAddrTemp= 1'b1; cif.ldCurrWordTemp = 1'b1; cif.hrq = 1'b1; end
        
	    state[iS2]: begin  cif.aen = 1'b1; cif.adstb = 1'b0; cif.checkReadWrite = 1'b1; cif.hrq = 1'b1; cif.checkWriteExtend = 1'b1; end
				

	    state[iS3]: begin cif.aen = 1'b1; cif.checkReadWrite = 1'b1; cif.hrq = 1'b1; end
		
	    state[iS4]: begin  cif.ldtempCurrAddr= 1'b1; cif.ldtempCurrWord = 1'b1; cif.validDACK = 1'b0;
			       cif.checkEOP = 1'b1; {cif.hrq, cif.aen} = 2'b00;
			end
					
    endcase
end
				 
endmodule		

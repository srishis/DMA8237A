// DMA Top module

module Dma8237aTop(dma_if.DUT dif, input logic CLK, RESET);


// DMA interface instantiation
DmaControlIf cif(CLK, RESET);

logic [5:0]  modeReg[4];
logic [7:0]  commandReg;
logic [7:0]  requestReg;
logic [7:0]  maskReg;

// DMA modules instantiation
// Datapath module
DmaDatapath D1(
		dp_if.DP, 
		cif, 
		.modeReg(modeReg), 
		.commandReg(commandReg),
		.requestReg(requestReg),
		.maskReg(maskReg)
);
	
	
// Timing and Control module
DmaTimingControl C1(
		     dif.TC, 
		     cif, 
		     .modeReg(modeReg), 
		     .commandReg(commandReg)
);

// Priority logic
DmaPriority P1(
		dif.PR, 
		.commandReg(commandReg),
		.requestReg(requestReg),
		.maskReg(maskReg)
);

endmodule

interface dmaRegIf(input logic CLK, RESET);

	logic [15:0] currAddrReg[0];
	logic [15:0] currAddrReg[1];
	logic [15:0] currAddrReg[2];
	logic [15:0] currAddrReg[3];
	logic [15:0] currWordReg[0];
	logic [15:0] currWordReg[1];
	logic [15:0] currWordReg[2];
	logic [15:0] currWordReg[3];
	logic [15:0] baseAddrReg[0];
	logic [15:0] baseAddrReg[1];
	logic [15:0] baseAddrReg[2];
	logic [15:0] baseAddrReg[3];
	logic [15:0] baseWordReg[0];
	logic [15:0] baseWordReg[1];
	logic [15:0] baseWordReg[2];
	logic [15:0] baseWordReg[3];
	logic [7:0]  modeReg[0];
	logic [7:0]  modeReg[1];
	logic [7:0]  modeReg[2];
	logic [7:0]  modeReg[3];
	logic [7:0]  commandReg;
	logic [7:0]  requestReg;
	logic [7:0]  maskReg;
	logic [7:0]  tempReg;
	logic [7:0]  statusReg;

endinterface
